`timescale 1ns / 1ps

module CSRRegs(
    input clk, rst,
    input[11:0] raddr, waddr,
    input[31:0] wdata,
    input csr_w,
    input[1:0] csr_wsc_mode,
    input[1:0] modifymip,
    input change,
    output[31:0] rdata,
    output sinterrupt,
    output[31:0] mstatus,
    output[31:0] mie
);

    reg[31:0] CSR [0:15];

    // Address mapping. The address is 12 bits, but only 4 bits are used in this module.
    wire raddr_valid = raddr[11:7] == 5'h6 && raddr[5:3] == 3'h0;
    wire[3:0] raddr_map = (raddr[6] << 3) + raddr[2:0];
    wire waddr_valid = waddr[11:7] == 5'h6 && waddr[5:3] == 3'h0;
    wire[3:0] waddr_map = (waddr[6] << 3) + waddr[2:0];

    assign mstatus = CSR[0];
    assign mie = CSR[4];
    assign sinterrupt = CSR[1][0];

    assign rdata = CSR[raddr_map];

    always@(posedge clk or posedge rst) begin
        if(rst) begin
			CSR[0] <= 32'h88;
			CSR[1] <= 0;
			CSR[2] <= 0;
			CSR[3] <= 0;
			CSR[4] <= 32'hfff;
			CSR[5] <= 0;
			CSR[6] <= 0;
			CSR[7] <= 0;
			CSR[8] <= 0;
			CSR[9] <= 0;
			CSR[10] <= 0;
			CSR[11] <= 0;
			CSR[12] <= 0;
			CSR[13] <= 0;
			CSR[14] <= 0;
			CSR[15] <= 0;
		end
        else if(csr_w || change) begin
            if(csr_w) begin
                case(csr_wsc_mode)
                    2'b01: CSR[waddr_map] = wdata;
                    2'b10: CSR[waddr_map] = CSR[waddr_map] | wdata;
                    2'b11: CSR[waddr_map] = CSR[waddr_map] & ~wdata;
                    default: CSR[waddr_map] = wdata;
                endcase
            end
            if(change) begin
                case(modifymip)
                    2'b00: begin
                        CSR[4] <= 32'hfff;
                    end
                    2'b01: begin
                        CSR[4] <= 32'hf7f;
                        if(~(|CSR[12])) CSR[12] <= CSR[9];
                        else begin
                            CSR[9] <= CSR[12];
                            CSR[12] <= 0;
                        end
                    end
                    2'b10: begin
                        CSR[4] <= 32'hf77;
                        if(~(|CSR[13])) CSR[13] <= CSR[9];
                        else begin
                            CSR[9] <= CSR[13];
                            CSR[13] <= 0;
                        end
                    end
                    2'b11: begin
                        CSR[4] <= 32'h777;
                        if(~(|CSR[14])) CSR[14] <= CSR[9];
                        else begin
                            CSR[9] <= CSR[14];
                            CSR[14] <= 0;
                        end
                    end
                endcase
            end
        end
    end
endmodule